library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity MyInstructionMemory is  
    port (
      Address : in std_logic_vector(31 downto 0);
      Instruction : out std_logic_vector(31 downto 0));
end entity MyInstructionMemory;

architecture Behavioral of MyInstructionMemory is
 type Memory is array (0 to 31) of std_logic_vector(31 downto 0);
 signal instructionMem : Memory := (
      "10001100000000110000000000000000", --1 lw $t3, 0($t0) -- t3 = 1
      "10001100000001000000000000000001", --2 lw $t4, 1($t0) -- t4 = 1
      "00000000011001000010000000000000", --3 add $t4, $t3, $t4
      "10101100000001000000000000000010", --4 sw $t4, 2($t0)
      "00000000011001000001100000000000", --5 add $t3, $t3, $t4
      "10101100000000110000000000000011", --6 sw $t3, 3($t0)
      "00000000011001000010000000000000", --7 add $t4, $t3, $t4
      "10101100000001000000000000000100", --8 sw $t4, 4($t0)
      "00000000011001000001100000000000", --9 add $t3, $t3, $t4
      "10101100000000110000000000000101", --10 sw $t3, 5($t0)
      "00000000011001000010000000000000", --11 add $t4, $t3, $t4
      "10101100000001000000000000000110", --12 sw $t4, 6($t0)
      "00000000011001000001100000000000", --13 add $t3, $t3, $t4
      "10101100000000110000000000000111", --14 sw $t3, 7($t0)         
      "00000000011001000010000000000000", --15 add $t4, $t3, $t4
      "10101100000001000000000000001000", --16 sw $t4, 8($t0) 
      "00000000011001000001100000000000", --17 add $t3, $t3, $t4
      "10101100000000110000000000001001", --18 sw $t3, 9($t0)
      "00000000011001000010000000000000", --19 add $t4, $t3, $t4
      "10101100000001000000000000001010", --20 sw $t4, 10($t0)
      "00000000000000000000000000000000", --21 Stall
      "00000000000000000000000000000000", --22 Stall
      "00000000000000000000000000000000", --23 Stall
      "00000000000000000000000000000000", --24 Stall
      "00000000000000000000000000000000", --25 Stall
      "00000000000000000000000000000000", --26 Stall	
      "00000000000000000000000000000000", --27 Stall
      "00000000000000000000000000000000", --28 Stall
      "00000000000000000000000000000000", --29 Stall	
      "00000000000000000000000000000000", --30 Stall
      "00000000000000000000000000000000", --31 Stall
      "00000000000000000000000000000000"); --32 Stall		

begin

 process(Address)
  begin
    report "Instruction Address = " & integer'image(to_integer(unsigned(Address)));
    Instruction <= instructionMem(to_integer(unsigned(Address)) / 4);
  end process;
           
end architecture Behavioral;



	

	

		
		





  



 

